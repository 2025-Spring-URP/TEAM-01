module ();
    initial begin
        $display("Hello, World!");
    end
endmodule